`timescale 1ns / 1ps
`include "define.svh"

import BasicTypes::*;
import PipelineTypes::*;

module Debug(
  DebugIF.Debug port
);

endmodule
