`timescale 1ns / 1ps
`include "define.svh"

module tracer(
  
);
endmodule
